LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY switch_2x2 IS
	PORT (
		X: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Y: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		V: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		C: OUT STD_LOGIC
	);
END switch_2x2;

ARCHITECTURE arch_switch_2x2 OF switch_2x2 IS
BEGIN
		U <= Y WHEN X(TO_INTEGER(UNSIGNED(S))) = '1' ELSE X;
		V <= X WHEN X(TO_INTEGER(UNSIGNED(S))) = '1' ELSE Y;
		C <= X(TO_INTEGER(UNSIGNED(S))) XNOR Y(TO_INTEGER(UNSIGNED(S)));
END ARCHITECTURE;
  